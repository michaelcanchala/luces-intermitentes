library verilog;
use verilog.vl_types.all;
entity rom_vlg_vec_tst is
end rom_vlg_vec_tst;
