library verilog;
use verilog.vl_types.all;
entity lucesintermitentes_vlg_check_tst is
    port(
        LD              : in     vl_logic;
        LI              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lucesintermitentes_vlg_check_tst;
