library verilog;
use verilog.vl_types.all;
entity lucesintermitentes_vlg_vec_tst is
end lucesintermitentes_vlg_vec_tst;
